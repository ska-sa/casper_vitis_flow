-- dsp_parameters.vhd 17. July 2018 by claus

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

LIBRARY UNISIM;
USE UNISIM.VComponents.all;

PACKAGE dsp_parameters IS

  SUBTYPE SHORT IS INTEGER RANGE 0 TO 1023;


  CONSTANT VERSION                      : STD_LOGIC_VECTOR(15 DOWNTO 0) := X"0000";

  CONSTANT HEADER_LAST_WORD_VALID_CONST : INTEGER  := 50;
--  CONSTANT HEADER_LAST_WORD_VALID_CONST : INTEGER  := 2;

  CONSTANT FRAGMENT1                    : INTEGER := 512 - HEADER_LAST_WORD_VALID_CONST * 8;
  CONSTANT FRAGMENT2                    : INTEGER := 512 - FRAGMENT1;

  CONSTANT TRUE                         : STD_LOGIC := '1';

END PACKAGE dsp_parameters;
